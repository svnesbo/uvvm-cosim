-- Todo
